`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/20/2025 08:58:18 PM
// Design Name: 
// Module Name: AddRound
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module AddRoundKey(

    input wire [127:0] state_in,
    input wire [127:0] round_key,
    output wire [127:0] state_out
    );
    
    assign state_out = state_in ^ round_key;
endmodule
